// program 1: 
`include "data_mem.sv"
`include "Top_level0.sv"
`include "new_fix2flt_tb.sv"

// program 2
/*
`include "data_mem.sv"
`include "flt2fix0.sv"
`include "flt2fix_tb.sv"
*/

// program 3
/*
`include "data_mem.sv"
`include "fltflt0_no_rnd.sv"
`include "fltflt_no_rnd_tb.sv"
*/

// `include "fltflt0_no_rnd.sv"
// `include "fltflt_no_rnd_tb.sv"